module xnor_test (a, b, out);
	input logic  a, b;
	output logic out;
endmodule