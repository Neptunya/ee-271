module pixel_selected (reset, left, right, row_select, current_pixel, next_pixel)


endmodule